// Assembly bytecode constants

`define NOP (32'h0000000)